library dot_matrix_sim;
package constants is
 
    constant clock_period : time := 0.25 ns; 
   
end package; 